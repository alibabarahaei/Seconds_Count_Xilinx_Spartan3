
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity clock_vhdl_module is
    Port ( clock : in  STD_LOGIC;
           out_1s : out  STD_LOGIC);
end clock_vhdl_module;

architecture Behavioral of clock_vhdl_module is

begin


end Behavioral;

